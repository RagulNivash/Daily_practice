`include "uvm_macros.svh"
import uvm_pkg::*;

class uart_config extends uvm_object;
  `uvm_object_utils(uart_config)

  function new(string name="uart_congif");
    super.new(name);
  endfunction

  uvm_active_passive_enum is_active=UVM_ACTIVE;

endclass


typedef enum bit[3:0] {rand_baud_1_stop=0,rand_length_1_stop=1, length5wp=2, length6wp=3, length7wp=4, length8wp=5, length5wop=6, length6wop=7, length7wop=8, length8wop=9, rand_baud_2_stop=11, rand_length_2_stop=12}oper_mode;

class transaction extends uvm_sequence_item;
  `uvm_object_utils(transaction)

rand oper mode op;
  logic tx_start, rx_start;
  logic rst;
  rand logic [16:0] baud;
  rand logic [7:0]tx_data;
  rand logic[3:0] length
  rand logic parity_type, parity_en;
  logic_stop2;
  logic t-done, rx_done, tx-err, rx_err;
  logic [7:0] rx_out;


  constraint baud_c{baud inside {4800, 9600, 14400, 19200, 38400, 57600};}
  constraint length_c {length inside {5,6,7,8};};

  function new(string name= "transaction");
    super.new(name);
  endfunction


endclass

////////////////////////////////////////////////////////////////////////////////////////////


class rand_baud extends uvm_sequence#(transaction);
  `uvm_object_utils(rand_baud)

  transaction tr;

  function new(string name="rand_baud");
    super.new(name);

  endfunction


  virtual task body();
    repeat(5)
      begin
        tr= transaction::type_ide::create("tr");
        start_item(tr);

      end


  endtask
      
    
